module prog(adres,out);

input [4:0] adres;
output [31:0] out;
reg [31:0] out;
 
reg [31:0] pmem [31:0];

always @(*)

begin
	out=pmem[adres];
end

initial
begin
 pmem[0]=32'b10000000010000000000000000000001;
 pmem[1]=32'b10000000100000000000000000000010;
 pmem[2]=32'b10000000110000000000000000000011;
 pmem[3]=32'b10000001000000000000000000000100;
 pmem[4]=32'b10000001010000000000000000000101;
 pmem[5]=32'b10000001100000000000000000000110;
 pmem[6]=32'b10000001110000000000000000000111;
 pmem[7]=32'b10000010000000000000000000001000;
 pmem[8]=32'b10000010010000000000000000001001;
 pmem[9]=32'b10000010100000000000000000001010;
pmem[10]=32'b10000010110000000000000000001011;
pmem[11]=32'b10000011000000000000000000001100;
pmem[12]=32'b10000011010000000000000000001101;
pmem[13]=32'b10000011100000000000000000001110;
pmem[14]=32'b10000011110000000000000000001111;
pmem[15]=32'b10000100000000000000000000010000;

pmem[16]=32'b00101000100000000000000101000010;
pmem[17]=32'b00101000110000000000000101100011;
pmem[18]=32'b00101001000000000000000110000100;
pmem[19]=32'b00101001010000000000000110100101;
pmem[20]=32'b00101001100000000000000111000110;
pmem[21]=32'b00101001110000000000000111100111;
pmem[22]=32'b00101010000000000000001000001000;


end
endmodule
