`include "mem.v"

//Deref is a module that performs load and store instructions and also passes the relevant raw values to the alu
module deref(opcode, rsrc1, rsrc2, enable, r );
endmodule
