module dot(gout,gl,al,gr);
	output gout;
	input gr,gl,al;
	assign gout = gl | (al & gr);
endmodule

module circle(gout,aout,gl,al,gr,ar);

	output gout,aout;
	input gl,al,gr,ar;
	assign gout = gl | (al & gr);
	assign aout = al & ar;

endmodule


module prefix(x,y,c,cout,s,clk);

	input[31:0]x,y;input c,clk;
	output[31:0]s;output cout;
	wire[31:0]p,g,a,l,p1,p2,p3,p4;
	wire[31:0]w1;
	wire [100:0]w2;
	wire [100:0]l1,l2,l3,l4,l5;

	assign p = x ^ y;
	assign g = x & y;
	assign a = g | p;
	assign w1[0]=c;

	dot d1(w1[1],g[0],a[0],c);
	
	circle c1(w2[1],w2[2],g[2],a[2],g[1],a[1]);
	circle c2(w2[3],w2[4],g[4],a[4],g[3],a[3]);
	circle c3(w2[5],w2[6],g[6],a[6],g[5],a[5]);
	circle c4(w2[7],w2[8],g[8],a[8],g[7],a[7]);
	circle c5(w2[9],w2[10],g[10],a[10],g[9],a[9]);
	circle c6(w2[11],w2[12],g[12],a[12],g[11],a[11]);
	circle c7(w2[13],w2[14],g[14],a[14],g[13],a[13]);
	circle c8(w2[15],w2[16],g[16],a[16],g[15],a[15]);
	circle c9(w2[17],w2[18],g[18],a[18],g[17],a[17]);
	circle c10(w2[19],w2[20],g[20],a[20],g[19],a[19]);
	circle c11(w2[21],w2[22],g[22],a[22],g[21],a[21]);
	circle c12(w2[23],w2[24],g[24],a[24],g[23],a[23]);
	circle c13(w2[25],w2[26],g[26],a[26],g[25],a[25]);
	circle c14(w2[27],w2[28],g[28],a[28],g[27],a[27]);
	circle c15(w2[29],w2[30],g[30],a[30],g[29],a[29]);

	dff f1(l1[0],clk,w1[0]);
	dff f2(l1[1],clk,w1[1]);
	dff f3(l1[2],clk,g[1]);
	dff f4(l1[3],clk,a[1]);
	dff f5(l1[4],clk,w2[1]);
	dff f6(l1[5],clk,w2[2]);
	dff f7(l1[6],clk,g[3]);
	dff f8(l1[7],clk,a[3]);
	dff f9(l1[8],clk,w2[3]);
	dff f10(l1[9],clk,w2[4]);
	dff f11(l1[10],clk,g[5]);
	dff f12(l1[11],clk,a[5]);
	dff f13(l1[12],clk,w2[5]);
	dff f14(l1[13],clk,w2[6]);
	dff f15(l1[14],clk,g[7]);
	dff f16(l1[15],clk,a[7]);
	dff f17(l1[16],clk,w2[7]);
	dff f18(l1[17],clk,w2[8]);
	dff f19(l1[18],clk,g[9]);
	dff f20(l1[19],clk,a[9]);
	dff f21(l1[20],clk,w2[9]);
	dff f22(l1[21],clk,w2[10]);
	dff f23(l1[22],clk,g[11]);
	dff f24(l1[23],clk,a[11]);
	dff f25(l1[24],clk,w2[11]);
	dff f26(l1[25],clk,w2[12]);
	dff f27(l1[26],clk,g[13]);
	dff f28(l1[27],clk,a[13]);
	dff f29(l1[28],clk,w2[13]);
	dff f30(l1[29],clk,w2[14]);
	dff f31(l1[30],clk,g[15]);
	dff f32(l1[31],clk,a[15]);
	dff f33(l1[32],clk,w2[15]);
	dff f34(l1[33],clk,w2[16]);
	dff f35(l1[34],clk,g[17]);
	dff f36(l1[35],clk,a[17]);
	dff f37(l1[36],clk,w2[17]);
	dff f38(l1[37],clk,w2[18]);
	dff f39(l1[38],clk,g[19]);
	dff f40(l1[39],clk,a[19]);
	dff f41(l1[40],clk,w2[19]);
	dff f42(l1[41],clk,w2[20]);
	dff f43(l1[42],clk,g[21]);
	dff f44(l1[43],clk,a[21]);
	dff f45(l1[44],clk,w2[21]);
	dff f46(l1[45],clk,w2[22]);
	dff f47(l1[46],clk,g[23]);
	dff f48(l1[47],clk,a[23]);
	dff f49(l1[48],clk,w2[23]);
	dff f50(l1[49],clk,w2[24]);
	dff f51(l1[50],clk,g[25]);
	dff f52(l1[51],clk,a[25]);
	dff f53(l1[52],clk,w2[25]);
	dff f54(l1[53],clk,w2[26]);
	dff f55(l1[54],clk,g[27]);
	dff f56(l1[55],clk,a[27]);
	dff f57(l1[56],clk,w2[27]);
	dff f58(l1[57],clk,w2[28]);
	dff f59(l1[58],clk,g[29]);
	dff f60(l1[59],clk,a[29]);
	dff f61(l1[60],clk,w2[29]);
	dff f62(l1[61],clk,w2[30]);
	dff f63(l1[62],clk,g[31]);
	dff f64(l1[63],clk,a[31]);


	dff f65(l[0],clk,p[0]);
	dff f66(l[1],clk,p[1]);
	dff f67(l[2],clk,p[2]);
	dff f68(l[3],clk,p[3]);
	dff f69(l[4],clk,p[4]);
	dff f70(l[5],clk,p[5]);
	dff f71(l[6],clk,p[6]);
	dff f72(l[7],clk,p[7]);
	dff f73(l[8],clk,p[8]);
	dff f74(l[9],clk,p[9]);
	dff f75(l[10],clk,p[10]);
	dff f76(l[11],clk,p[11]);
	dff f77(l[12],clk,p[12]);
	dff f78(l[13],clk,p[13]);
	dff f79(l[14],clk,p[14]);
	dff f80(l[15],clk,p[15]);
	dff f81(l[16],clk,p[16]);
	dff f82(l[17],clk,p[17]);
	dff f83(l[18],clk,p[18]);
	dff f84(l[19],clk,p[19]);
	dff f85(l[20],clk,p[20]);
	dff f86(l[21],clk,p[21]);
	dff f87(l[22],clk,p[22]);
	dff f88(l[23],clk,p[23]);
	dff f89(l[24],clk,p[24]);
	dff f90(l[25],clk,p[25]);
	dff f91(l[26],clk,p[26]);
	dff f92(l[27],clk,p[27]);
	dff f93(l[28],clk,p[28]);
	dff f94(l[29],clk,p[29]);
	dff f95(l[30],clk,p[30]);
	dff f96(l[31],clk,p[31]);

	dot d2(w1[2],l1[2],l1[3],l1[1]);
	dot d3(w1[3],l1[4],l1[5],l1[1]);

	circle c16(w2[31],w2[32],l1[10],l1[11],l1[8],l1[9]);
	circle c17(w2[33],w2[34],l1[12],l1[13],l1[8],l1[9]);
	circle c18(w2[35],w2[36],l1[18],l1[19],l1[16],l1[17]);
	circle c19(w2[37],w2[38],l1[20],l1[21],l1[16],l1[17]);
	circle c20(w2[39],w2[40],l1[26],l1[27],l1[24],l1[25]);
	circle c21(w2[41],w2[42],l1[28],l1[29],l1[24],l1[25]);
	circle c22(w2[43],w2[44],l1[34],l1[35],l1[32],l1[33]);
	circle c23(w2[45],w2[46],l1[36],l1[37],l1[32],l1[33]);
	circle c24(w2[47],w2[48],l1[42],l1[43],l1[40],l1[41]);
	circle c25(w2[49],w2[50],l1[44],l1[45],l1[40],l1[41]);
	circle c26(w2[51],w2[52],l1[50],l1[51],l1[48],l1[49]);
	circle c27(w2[53],w2[54],l1[52],l1[53],l1[48],l1[49]);
	circle c28(w2[55],w2[56],l1[58],l1[59],l1[56],l1[57]);
	circle c29(w2[57],w2[58],l1[60],l1[61],l1[56],l1[57]);

	dff b1(l2[0],clk,l1[0]);
	dff b2(l2[1],clk,l1[1]);
	dff b3(l2[2],clk,w1[2]);
	dff b4(l2[3],clk,w1[3]);
	dff b5(l2[4],clk,l1[6]);
	dff b6(l2[5],clk,l1[7]);
	dff b7(l2[6],clk,l1[8]);
	dff b8(l2[7],clk,l1[9]);
	dff b9(l2[8],clk,w2[31]);
	dff b10(l2[9],clk,w2[32]);
	dff b11(l2[10],clk,w2[33]);
	dff b12(l2[11],clk,w2[34]);
	dff b13(l2[12],clk,l1[14]);
	dff b14(l2[13],clk,l1[15]);
	dff b15(l2[14],clk,l1[16]);
	dff b16(l2[15],clk,l1[17]);
	dff b17(l2[16],clk,w2[35]);
	dff b18(l2[17],clk,w2[36]);
	dff b19(l2[18],clk,w2[37]);
	dff b20(l2[19],clk,w2[38]);
	dff b21(l2[20],clk,l1[22]);
	dff b22(l2[21],clk,l1[23]);
	dff b23(l2[22],clk,l1[24]);
	dff b24(l2[23],clk,l1[25]);
	dff b25(l2[24],clk,w2[39]);
	dff b26(l2[25],clk,w2[40]);
	dff b27(l2[26],clk,w2[41]);
	dff b28(l2[27],clk,w2[42]);
	dff b29(l2[28],clk,l1[30]);
	dff b30(l2[29],clk,l1[31]);
	dff b31(l2[30],clk,l1[32]);
	dff b32(l2[31],clk,l1[33]);
	dff b33(l2[32],clk,w2[43]);
	dff b34(l2[33],clk,w2[44]);
	dff b35(l2[34],clk,w2[45]);
	dff b36(l2[35],clk,w2[46]);
	dff b37(l2[36],clk,l1[38]);
	dff b38(l2[37],clk,l1[39]);
	dff b39(l2[38],clk,l1[40]);
	dff b40(l2[39],clk,l1[41]);
	dff b41(l2[40],clk,w2[47]);
	dff b42(l2[41],clk,w2[48]);
	dff b43(l2[42],clk,w2[49]);
	dff b44(l2[43],clk,w2[50]);
	dff b45(l2[44],clk,l1[46]);
	dff b46(l2[45],clk,l1[47]);
	dff b47(l2[46],clk,l1[48]);
	dff b48(l2[47],clk,l1[49]);
	dff b49(l2[48],clk,w2[51]);
	dff b50(l2[49],clk,w2[52]);
	dff b51(l2[50],clk,w2[53]);
	dff b52(l2[51],clk,w2[54]);
	dff b53(l2[52],clk,l1[54]);
	dff b54(l2[53],clk,l1[55]);
	dff b55(l2[54],clk,l1[56]);
	dff b56(l2[55],clk,l1[57]);
	dff b57(l2[56],clk,w2[55]);
	dff b58(l2[57],clk,w2[56]);
	dff b59(l2[58],clk,w2[57]);
	dff b60(l2[59],clk,w2[58]);
	dff b61(l2[60],clk,l1[62]);
	dff b62(l2[61],clk,l1[63]);

	dff b65 (p1[0],clk,l[0]);
	dff b66 (p1[1],clk,l[1]);
	dff b67 (p1[2],clk,l[2]);
	dff b68 (p1[3],clk,l[3]);
	dff b69 (p1[4],clk,l[4]);
	dff b70 (p1[5],clk,l[5]);
	dff b71 (p1[6],clk,l[6]);
	dff b72 (p1[7],clk,l[7]);
	dff b73 (p1[8],clk,l[8]);
	dff b74 (p1[9],clk,l[9]);
	dff b75 (p1[10],clk,l[10]);
	dff b76 (p1[11],clk,l[11]);
	dff b77 (p1[12],clk,l[12]);
	dff b78 (p1[13],clk,l[13]);
	dff b79 (p1[14],clk,l[14]);
	dff b80 (p1[15],clk,l[15]);
	dff b81 (p1[16],clk,l[16]);
	dff b82 (p1[17],clk,l[17]);
	dff b83 (p1[18],clk,l[18]);
	dff b84 (p1[19],clk,l[19]);
	dff b85 (p1[20],clk,l[20]);
	dff b86 (p1[21],clk,l[21]);
	dff b87 (p1[22],clk,l[22]);
	dff b88 (p1[23],clk,l[23]);
	dff b89 (p1[24],clk,l[24]);
	dff b90 (p1[25],clk,l[25]);
	dff b91 (p1[26],clk,l[26]);
	dff b92 (p1[27],clk,l[27]);
	dff b93 (p1[28],clk,l[28]);
	dff b94 (p1[29],clk,l[29]);
	dff b95 (p1[30],clk,l[30]);
	dff b96 (p1[31],clk,l[31]);

	dot d4(w1[4],l2[4],l2[5],l2[3]);
	dot d5(w1[5],l2[6],l2[7],l2[3]);
	dot d6(w1[6],l2[8],l2[9],l2[3]);
	dot d7(w1[7],l2[10],l2[11],l2[3]);
	
	circle c30(w2[59],w2[60],l2[20],l2[21],l2[18],l2[19]);
	circle c31(w2[61],w2[62],l2[22],l2[23],l2[18],l2[19]);
	circle c32(w2[63],w2[64],l2[24],l2[25],l2[18],l2[19]);
	circle c33(w2[65],w2[66],l2[26],l2[27],l2[18],l2[19]);
	circle c34(w2[67],w2[68],l2[36],l2[37],l2[34],l2[35]);
	circle c35(w2[69],w2[70],l2[38],l2[39],l2[34],l2[35]);
	circle c36(w2[71],w2[72],l2[40],l2[41],l2[34],l2[35]);
	circle c37(w2[73],w2[74],l2[42],l2[43],l2[34],l2[35]);
	circle c38(w2[75],w2[76],l2[52],l2[53],l2[50],l2[51]);
	circle c39(w2[77],w2[78],l2[54],l2[55],l2[50],l2[51]);
	circle c40(w2[79],w2[80],l2[56],l2[57],l2[50],l2[51]);
	circle c41(w2[81],w2[82],l2[58],l2[59],l2[50],l2[51]);

	dff m1(l3[0],clk,l2[0]);
	dff m2(l3[1],clk,l2[1]);
	dff m3(l3[2],clk,l2[2]);
	dff m4(l3[3],clk,l2[3]);
	dff m5(l3[4],clk,w1[4]);
	dff m6(l3[5],clk,w1[5]);
	dff m7(l3[6],clk,w1[6]);
	dff m8(l3[7],clk,w1[7]);
	dff m9(l3[8],clk,l2[12]);
	dff m10(l3[9],clk,l2[13]);
	dff m11(l3[10],clk,l2[14]);
	dff m12(l3[11],clk,l2[15]);
	dff m13(l3[12],clk,l2[16]);
	dff m14(l3[13],clk,l2[17]);
	dff m15(l3[14],clk,l2[18]);
	dff m16(l3[15],clk,l2[19]);
	dff m17(l3[16],clk,w2[59]);
	dff m18(l3[17],clk,w2[60]);
	dff m19(l3[18],clk,w2[61]);
	dff m20(l3[19],clk,w2[62]);
	dff m21(l3[20],clk,w2[63]);
	dff m22(l3[21],clk,w2[64]);
	dff m23(l3[22],clk,w2[65]);
	dff m24(l3[23],clk,w2[66]);
	dff m25(l3[24],clk,l2[28]);
	dff m26(l3[25],clk,l2[29]);
	dff m27(l3[26],clk,l2[30]);
	dff m28(l3[27],clk,l2[31]);
	dff m29(l3[28],clk,l2[32]);
	dff m30(l3[29],clk,l2[33]);
	dff m31(l3[30],clk,l2[34]);
	dff m32(l3[31],clk,l2[35]);
	dff m33(l3[32],clk,w2[67]);
	dff m34(l3[33],clk,w2[68]);
	dff m35(l3[34],clk,w2[69]);
	dff m36(l3[35],clk,w2[70]);
	dff m37(l3[36],clk,w2[71]);
	dff m38(l3[37],clk,w2[72]);
	dff m39(l3[38],clk,w2[73]);
	dff m40(l3[39],clk,w2[74]);
	dff m41(l3[40],clk,l2[44]);
	dff m42(l3[41],clk,l2[45]);
	dff m43(l3[42],clk,l2[46]);
	dff m44(l3[43],clk,l2[47]);
	dff m45(l3[44],clk,l2[48]);
	dff m46(l3[45],clk,l2[49]);
	dff m47(l3[46],clk,l2[50]);
	dff m48(l3[47],clk,l2[51]);
	dff m49(l3[48],clk,w2[75]);
	dff m50(l3[49],clk,w2[76]);
	dff m51(l3[50],clk,w2[77]);
	dff m52(l3[51],clk,w2[78]);
	dff m53(l3[52],clk,w2[79]);
	dff m54(l3[53],clk,w2[80]);
	dff m55(l3[54],clk,w2[81]);
	dff m56(l3[56],clk,w2[82]);
	dff m57(l3[56],clk,l2[60]);
	dff m58(l3[57],clk,l2[61]);

	dff m65 (p2[0],clk,p1[0]);
	dff m66 (p2[1],clk,p1[1]);
	dff m67 (p2[2],clk,p1[2]);
	dff m68 (p2[3],clk,p1[3]);
	dff m69 (p2[4],clk,p1[4]);
	dff m70 (p2[5],clk,p1[5]);
	dff m71 (p2[6],clk,p1[6]);
	dff m72 (p2[7],clk,p1[7]);
	dff m73 (p2[8],clk,p1[8]);
	dff m74 (p2[9],clk,p1[9]);
	dff m75 (p2[10],clk,p1[10]);
	dff m76 (p2[11],clk,p1[11]);
	dff m77 (p2[12],clk,p1[12]);
	dff m78 (p2[13],clk,p1[13]);
	dff m79 (p2[14],clk,p1[14]);
	dff m80 (p2[15],clk,p1[15]);
	dff m81 (p2[16],clk,p1[16]);
	dff m82 (p2[17],clk,p1[17]);
	dff m83 (p2[18],clk,p1[18]);
	dff m84 (p2[19],clk,p1[19]);
	dff m85 (p2[20],clk,p1[20]);
	dff m86 (p2[21],clk,p1[21]);
	dff m87 (p2[22],clk,p1[22]);
	dff m88 (p2[23],clk,p1[23]);
	dff m89 (p2[24],clk,p1[24]);
	dff m90 (p2[25],clk,p1[25]);
	dff m91 (p2[26],clk,p1[26]);
	dff m92 (p2[27],clk,p1[27]);
	dff m93 (p2[28],clk,p1[28]);
	dff m94 (p2[29],clk,p1[29]);
	dff m95 (p2[30],clk,p1[30]);
	dff m96 (p2[31],clk,p1[31]);

	dot d8(w1[8],l3[8],l3[9],l3[7]);
	dot d9(w1[9],l3[10],l3[11],l3[7]);
	dot d10(w1[10],l3[12],l3[13],l3[7]);
	dot d11(w1[11],l3[14],l3[15],l3[7]);
	dot d12(w1[12],l3[16],l3[17],l3[7]);
	dot d13(w1[13],l3[18],l3[19],l3[7]);
	dot d14(w1[14],l3[20],l3[21],l3[7]);
	dot d15(w1[15],l3[22],l3[23],l3[7]);
	circle c42(w2[83],w2[84],l3[40],l3[41],l3[38],l3[39]);
	circle c43(w2[85],w2[86],l3[42],l3[43],l3[38],l3[39]);
	circle c44(w2[87],w2[88],l3[44],l3[45],l3[38],l3[39]);
	circle c45(w2[89],w2[90],l3[46],l3[47],l3[38],l3[39]);
	circle c46(w2[91],w2[92],l3[48],l3[49],l3[38],l3[39]);
	circle c47(w2[93],w2[94],l3[50],l3[51],l3[38],l3[39]);
	circle c48(w2[95],w2[96],l3[52],l3[53],l3[38],l3[39]);
	circle c49(w2[97],w2[98],l3[54],l3[55],l3[38],l3[39]);

	dff z1(l4[0],clk,l3[0]);
	dff z2(l4[1],clk,l3[1]);
	dff z3(l4[2],clk,l3[2]);
	dff z4(l4[3],clk,l3[3]);
	dff z5(l4[4],clk,l3[4]);
	dff z6(l4[5],clk,l3[5]);
	dff z7(l4[6],clk,l3[6]);
	dff z8(l4[7],clk,l3[7]);
	dff z9(l4[8],clk,w1[8]);
	dff z10(l4[9],clk,w1[9]);
	dff z11(l4[10],clk,w1[10]);
	dff z12(l4[11],clk,w1[11]);
	dff z13(l4[12],clk,w1[12]);
	dff z14(l4[13],clk,w1[13]);
	dff z15(l4[14],clk,w1[14]);
	dff z16(l4[15],clk,w1[15]);
	dff z17(l4[16],clk,l3[24]);
	dff z18(l4[17],clk,l3[25]);
	dff z19(l4[18],clk,l3[26]);
	dff z20(l4[19],clk,l3[27]);
	dff z21(l4[20],clk,l3[28]);
	dff z22(l4[21],clk,l3[29]);
	dff z23(l4[22],clk,l3[30]);
	dff z24(l4[23],clk,l3[31]);
	dff z25(l4[24],clk,l3[32]);
	dff z26(l4[25],clk,l3[33]);
	dff z27(l4[26],clk,l3[34]);
	dff z28(l4[27],clk,l3[35]);
	dff z29(l4[28],clk,l3[36]);
	dff z30(l4[29],clk,l3[37]);
	dff z31(l4[30],clk,l3[38]);
	dff z32(l4[31],clk,l3[39]);
	dff z33(l4[32],clk,w2[83]);
	dff z34(l4[33],clk,w2[84]);
	dff z35(l4[34],clk,w2[85]);
	dff z36(l4[35],clk,w2[86]);
	dff z37(l4[36],clk,w2[87]);
	dff z38(l4[37],clk,w2[88]);
	dff z39(l4[38],clk,w2[89]);
	dff z40(l4[39],clk,w2[90]);
	dff z41(l4[40],clk,w2[91]);
	dff z42(l4[41],clk,w2[92]);
	dff z43(l4[42],clk,w2[93]);
	dff z44(l4[43],clk,w2[94]);
	dff z45(l4[44],clk,w2[95]);
	dff z46(l4[45],clk,w2[96]);
	dff z47(l4[46],clk,w2[97]);
	dff z48(l4[47],clk,w2[98]);
	dff z49(l4[48],clk,l3[56]);
	dff z50(l4[49],clk,l3[57]);

	dff n65 (p3[0],clk,p2[0]);
	dff n66 (p3[1],clk,p2[1]);
	dff n67 (p3[2],clk,p2[2]);
	dff n68 (p3[3],clk,p2[3]);
	dff n69 (p3[4],clk,p2[4]);
	dff n70 (p3[5],clk,p2[5]);
	dff n71 (p3[6],clk,p2[6]);
	dff n72 (p3[7],clk,p2[7]);
	dff n73 (p3[8],clk,p2[8]);
	dff n74 (p3[9],clk,p2[9]);
	dff n75 (p3[10],clk,p2[10]);
	dff n76 (p3[11],clk,p2[11]);
	dff n77 (p3[12],clk,p2[12]);
	dff n78 (p3[13],clk,p2[13]);
	dff n79 (p3[14],clk,p2[14]);
	dff n80 (p3[15],clk,p2[15]);
	dff n81 (p3[16],clk,p2[16]);
	dff n82 (p3[17],clk,p2[17]);
	dff n83 (p3[18],clk,p2[18]);
	dff n84 (p3[19],clk,p2[19]);
	dff n85 (p3[20],clk,p2[20]);
	dff n86 (p3[21],clk,p2[21]);
	dff n87 (p3[22],clk,p2[22]);
	dff n88 (p3[23],clk,p2[23]);
	dff n89 (p3[24],clk,p2[24]);
	dff n90 (p3[25],clk,p2[25]);
	dff n91 (p3[26],clk,p2[26]);
	dff n92 (p3[27],clk,p2[27]);
	dff n93 (p3[28],clk,p2[28]);
	dff n94 (p3[29],clk,p2[29]);
	dff n95 (p3[30],clk,p2[30]);
	dff n96 (p3[31],clk,p2[31]);

	dot d16(w1[16],l4[16],l4[17],l4[15]);
	dot d17(w1[17],l4[18],l4[19],l4[15]);
	dot d18(w1[18],l4[20],l4[21],l4[15]);
	dot d19(w1[19],l4[22],l4[23],l4[15]);
	dot d20(w1[20],l4[24],l4[25],l4[15]);
	dot d21(w1[21],l4[26],l4[27],l4[15]);
	dot d22(w1[22],l4[28],l4[29],l4[15]);
	dot d23(w1[23],l4[30],l4[31],l4[15]);
	dot d24(w1[24],l4[32],l4[33],l4[15]);
	dot d25(w1[25],l4[34],l4[35],l4[15]);
	dot d26(w1[26],l4[36],l4[37],l4[15]);
	dot d27(w1[27],l4[38],l4[39],l4[15]);
	dot d28(w1[28],l4[40],l4[41],l4[15]);
	dot d29(w1[29],l4[42],l4[43],l4[15]);
	dot d30(w1[30],l4[44],l4[45],l4[15]);
	dot d31(w1[31],l4[46],l4[47],l4[15]);

	dff q1(l5[0],clk,l4[0]);
	dff q2(l5[1],clk,l4[1]);
	dff q3(l5[2],clk,l4[2]);
	dff q4(l5[3],clk,l4[3]);
	dff q5(l5[4],clk,l4[4]);
	dff q6(l5[5],clk,l4[5]);
	dff q7(l5[6],clk,l4[6]);
	dff q8(l5[7],clk,l4[7]);
	dff q9(l5[8],clk,l4[8]);
	dff q10(l5[9],clk,l4[9]);
	dff q11(l5[10],clk,l4[10]);
	dff q12(l5[11],clk,l4[11]);
	dff q13(l5[12],clk,l4[12]);
	dff q14(l5[13],clk,l4[13]);
	dff q15(l5[14],clk,l4[14]);
	dff q16(l5[15],clk,l4[15]);
	dff q17(l5[16],clk,w1[16]);
	dff q18(l5[17],clk,w1[17]);
	dff q19(l5[18],clk,w1[18]);
	dff q20(l5[19],clk,w1[19]);
	dff q21(l5[20],clk,w1[20]);
	dff q22(l5[21],clk,w1[21]);
	dff q23(l5[22],clk,w1[22]);
	dff q24(l5[23],clk,w1[23]);
	dff q25(l5[24],clk,w1[24]);
	dff q26(l5[25],clk,w1[25]);
	dff q27(l5[26],clk,w1[26]);
	dff q28(l5[27],clk,w1[27]);
	dff q29(l5[28],clk,w1[28]);
	dff q30(l5[29],clk,w1[29]);
	dff q31(l5[30],clk,w1[30]);
	dff q32(l5[31],clk,w1[31]);
	dff q33(l5[32],clk,l4[48]);
	dff q34(l5[33],clk,l4[49]);

	dff z65 (p4[0],clk,p3[0]);
	dff z66 (p4[1],clk,p3[1]);
	dff z67 (p4[2],clk,p3[2]);
	dff z68 (p4[3],clk,p3[3]);
	dff z69 (p4[4],clk,p3[4]);
	dff z70 (p4[5],clk,p3[5]);
	dff z71 (p4[6],clk,p3[6]);
	dff z72 (p4[7],clk,p3[7]);
	dff z73 (p4[8],clk,p3[8]);
	dff z74 (p4[9],clk,p3[9]);
	dff z75 (p4[10],clk,p3[10]);
	dff z76 (p4[11],clk,p3[11]);
	dff z77 (p4[12],clk,p3[12]);
	dff z78 (p4[13],clk,p3[13]);
	dff z79 (p4[14],clk,p3[14]);
	dff z80 (p4[15],clk,p3[15]);
	dff z81 (p4[16],clk,p3[16]);
	dff z82 (p4[17],clk,p3[17]);
	dff z83 (p4[18],clk,p3[18]);
	dff z84 (p4[19],clk,p3[19]);
	dff z85 (p4[20],clk,p3[20]);
	dff z86 (p4[21],clk,p3[21]);
	dff z87 (p4[22],clk,p3[22]);
	dff z88 (p4[23],clk,p3[23]);
	dff z89 (p4[24],clk,p3[24]);
	dff z90 (p4[25],clk,p3[25]);
	dff z91 (p4[26],clk,p3[26]);
	dff z92 (p4[27],clk,p3[27]);
	dff z93 (p4[28],clk,p3[28]);
	dff z94 (p4[29],clk,p3[29]);
	dff z95 (p4[30],clk,p3[30]);
	dff z96 (p4[31],clk,p3[31]);

	dot d32(cout,l5[32],l5[33],l5[31]);
	assign s = p4[31:0] ^ l5[31:0];

endmodule

