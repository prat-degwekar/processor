`include "fpa_adder.v"

module fpa_addertb();
	reg [31:0]a,b;
	reg  clk,inp_op;
	wire [31:0]out;

	fpa_adder f0(a,b,clk,inp_op,out);
	/*
	initial
	begin
	$monitor(" \t a: %b b:%b  out=%b\t",a,b,out);
	end
	*/
	initial
	begin
	    //$dumpfile("test.vcd");
	    //$dumpvars;
	    $monitor("a = %d , b = %d , inp_op = %b , out = %d\n",a , b , inp_op , out);
	end

	always begin

		#150

		$finish;

	end

	initial	begin
		clk=0;

		a=32'b01000000110111111010110001110001;    //6.9898     129
		b=32'b01000100011101101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=0;

		/*#10

		a=32'b11000000110111111010110010110001;    //6.9898     129
		b=32'b11000100011101101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=1;

		#10

		a=32'b11000000110111111010110001110001;    //6.9898     129
		b=32'b01000110011101101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=1;

		#10

		a=32'b01011000110111111010110001110001;    //6.9898     129
		b=32'b11000100011101101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=0;

		#10

		b=32'b01000000110111111010110001110001;    //6.9898     129
		a=32'b01011100011101101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=1;

		#10

		b=32'b11000000111111111010110001110001;    //6.9898     129
		a=32'b11000100011101101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=1;

		#10

		b=32'b11010000110111111010110001110001;    //6.9898     129
		a=32'b01000100011111101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=0;

		#10

		b=32'b01000000110111111010110001110001;    //6.9898     129
		a=32'b11001001011101101011100110010110;     //986.8998  136    //6.9898+986.8998

		inp_op=1;*/

	end
	
	 always begin
	 	#5
	 		clk = ~clk; // Toggle clock every 5 ticks
	 end
endmodule
