module pgen(a,b,c);

    input [31:0]a;
    input b;
    output [31:0]c;

    assign c[0]=a[0]&b;
    assign c[1]=a[1]&b;
    assign c[2]=a[2]&b;
    assign c[3]=a[3]&b;
    assign c[4]=a[4]&b;
    assign c[5]=a[5]&b;
    assign c[6]=a[6]&b;
    assign c[7]=a[7]&b;
    assign c[8]=a[8]&b;
    assign c[9]=a[9]&b;
    assign c[10]=a[10]&b;
    assign c[11]=a[11]&b;
    assign c[12]=a[12]&b;
    assign c[13]=a[13]&b;
    assign c[14]=a[14]&b;
    assign c[15]=a[15]&b;
    assign c[16]=a[16]&b;
    assign c[17]=a[17]&b;
    assign c[18]=a[18]&b;
    assign c[19]=a[19]&b;
    assign c[20]=a[20]&b;
    assign c[21]=a[21]&b;
    assign c[22]=a[22]&b;
    assign c[23]=a[23]&b;
    assign c[24]=a[24]&b;
    assign c[25]=a[25]&b;
    assign c[26]=a[26]&b;
    assign c[27]=a[27]&b;
    assign c[28]=a[28]&b;
    assign c[29]=a[29]&b;
    assign c[30]=a[30]&b;
    assign c[31]=a[31]&b;

endmodule
